`timescale 1ns / 1ps
module bcd7_ext();

endmodule